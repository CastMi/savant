architecture imp of andport is

begin
f <= a and b;
end architecture imp;

