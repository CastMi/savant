library ieee;
use ieee.std_logic_1164.all;

entity andport is
 port (
   signal a : in bit;
   signal b : in bit;
   signal f : out bit);
end entity andport;

