--
-- Copyright (c) 2015 Michele Castellana (michele.castellana@mail.polimi.it)
--
--    This source code is free software; you can redistribute it
--    and/or modify it in source code form under the terms of the GNU
--    General Public License as published by the Free Software
--    Foundation; either version 2 of the License, or (at your option)
--    any later version.
--
--    This program is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--
--    You should have received a copy of the GNU General Public License
--    along with this program; if not, write to the Free Software
--    Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA.
--

-- library declaration
library IEEE;
use IEEE.std_logic_1164.all;

-- entity
entity AndPort is Port (
	A, B : in bit;
	F  	 : out bit
	);
end AndPort;

-- architecture
architecture imp of AndPort is
	begin
		F <= A and B;
end imp;
